library verilog;
use verilog.vl_types.all;
entity upcount_vlg_vec_tst is
end upcount_vlg_vec_tst;
