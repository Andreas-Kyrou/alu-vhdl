library verilog;
use verilog.vl_types.all;
entity Project3_vlg_vec_tst is
end Project3_vlg_vec_tst;
